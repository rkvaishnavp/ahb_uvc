typedef class uvm_sequencer#(ahb_tx) ahb_sqr;