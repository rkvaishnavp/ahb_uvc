typedef uvm_sequencer#(ahb_tx) ahb_sqr;
